library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

-- Alpha-max-beta-min approximation: |Z| ≈ max + 0.375*min
-- Avoids CORDIC/sqrt, <4% error worst case

entity magnitude_calc is
    Generic (
        DATA_WIDTH : integer := 16;
        OUT_WIDTH  : integer := 17
    );
    Port (
        aclk          : in  STD_LOGIC;
        aresetn       : in  STD_LOGIC;
        s_axis_tdata  : in  STD_LOGIC_VECTOR(2*DATA_WIDTH-1 downto 0);
        s_axis_tvalid : in  STD_LOGIC;
        s_axis_tready : out STD_LOGIC;
        s_axis_tlast  : in  STD_LOGIC;
        m_axis_tdata  : out STD_LOGIC_VECTOR(OUT_WIDTH-1 downto 0);
        m_axis_tvalid : out STD_LOGIC;
        m_axis_tready : in  STD_LOGIC;
        m_axis_tlast  : out STD_LOGIC
    );
end magnitude_calc;

architecture Behavioral of magnitude_calc is

    signal s1_max, s1_min : unsigned(DATA_WIDTH-1 downto 0) := (others => '0');
    signal s1_valid       : std_logic := '0';
    signal s1_last        : std_logic := '0';
    
    signal s2_mag   : unsigned(OUT_WIDTH-1 downto 0) := (others => '0');
    signal s2_valid : std_logic := '0';
    signal s2_last  : std_logic := '0';
    
    signal pipe_enable : std_logic;

begin

    pipe_enable <= m_axis_tready or (not s2_valid);
    s_axis_tready <= pipe_enable;

    stage1_proc: process(aclk)
        variable i_signed, q_signed : signed(DATA_WIDTH-1 downto 0);
        variable abs_i, abs_q       : unsigned(DATA_WIDTH-1 downto 0);
    begin
        if rising_edge(aclk) then
            if aresetn = '0' then
                s1_max   <= (others => '0');
                s1_min   <= (others => '0');
                s1_valid <= '0';
                s1_last  <= '0';
            elsif pipe_enable = '1' then
                if s_axis_tvalid = '1' then
                    i_signed := signed(s_axis_tdata(DATA_WIDTH-1 downto 0));
                    q_signed := signed(s_axis_tdata(2*DATA_WIDTH-1 downto DATA_WIDTH));
                    
                    if i_signed(DATA_WIDTH-1) = '1' then
                        abs_i := unsigned(-i_signed);
                    else
                        abs_i := unsigned(i_signed);
                    end if;
                    
                    if q_signed(DATA_WIDTH-1) = '1' then
                        abs_q := unsigned(-q_signed);
                    else
                        abs_q := unsigned(q_signed);
                    end if;
                    
                    if abs_i >= abs_q then
                        s1_max <= abs_i;
                        s1_min <= abs_q;
                    else
                        s1_max <= abs_q;
                        s1_min <= abs_i;
                    end if;
                    
                    s1_valid <= '1';
                    s1_last  <= s_axis_tlast;
                else
                    s1_valid <= '0';
                    s1_last  <= '0';
                end if;
            end if;
        end if;
    end process;

    -- 0.375 = 1/4 + 1/8 = (min >> 2) + (min >> 3)
    stage2_proc: process(aclk)
        variable max_ext, min_div4, min_div8 : unsigned(OUT_WIDTH-1 downto 0);
    begin
        if rising_edge(aclk) then
            if aresetn = '0' then
                s2_mag   <= (others => '0');
                s2_valid <= '0';
                s2_last  <= '0';
            elsif pipe_enable = '1' then
                if s1_valid = '1' then
                    max_ext  := resize(s1_max, OUT_WIDTH);
                    min_div4 := resize(s1_min(DATA_WIDTH-1 downto 2), OUT_WIDTH);
                    min_div8 := resize(s1_min(DATA_WIDTH-1 downto 3), OUT_WIDTH);
                    s2_mag   <= max_ext + min_div4 + min_div8;
                    s2_valid <= '1';
                    s2_last  <= s1_last;
                else
                    s2_valid <= '0';
                    s2_last  <= '0';
                end if;
            end if;
        end if;
    end process;

    m_axis_tdata  <= std_logic_vector(s2_mag);
    m_axis_tvalid <= s2_valid;
    m_axis_tlast  <= s2_last;

end Behavioral;