library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.ALL;
use std.textio.all;
use IEEE.std_logic_textio.all;

-- =============================================================================
-- Testbench: Radar Core v3/v4 Verification (Optimized - No Magic Waits)
-- =============================================================================

entity tb_radar_core is
end tb_radar_core;

architecture Behavioral of tb_radar_core is

    component radar_core_v3 is
        Generic (
            N_RANGE   : integer := 1024;
            N_DOPPLER : integer := 128
        );
        Port (
            aclk            : in  STD_LOGIC;
            aresetn         : in  STD_LOGIC;
            s_axis_tdata    : in  STD_LOGIC_VECTOR(31 downto 0);
            s_axis_tvalid   : in  STD_LOGIC;
            s_axis_tlast    : in  STD_LOGIC;
            s_axis_tready   : out STD_LOGIC;
            m_axis_tdata    : out STD_LOGIC_VECTOR(16 downto 0);
            m_axis_tvalid   : out STD_LOGIC;
            m_axis_tlast    : out STD_LOGIC;
            m_axis_tready   : in  STD_LOGIC;
            rdm_range_bin   : out STD_LOGIC_VECTOR(9 downto 0);
            rdm_doppler_bin : out STD_LOGIC_VECTOR(6 downto 0);
            status_range_fft_done   : out STD_LOGIC;
            status_doppler_fft_done : out STD_LOGIC;
            status_frame_complete   : out STD_LOGIC;
            status_overflow         : out STD_LOGIC
        );
    end component;

    -- =========================================================================
    -- Test Parameters
    -- =========================================================================
    constant N_RANGE    : integer := 1024;
    constant N_DOPPLER  : integer := 128;
    constant CLK_PERIOD : time := 10 ns;
    
    -- Target parameters
    constant TARGET_1_RANGE   : integer := 100;
    constant TARGET_1_DOPPLER : real := 5.0;
    constant TARGET_1_AMP     : real := 8000.0;
    
    constant TARGET_2_RANGE   : integer := 500;
    constant TARGET_2_DOPPLER : real := -10.0;
    constant TARGET_2_AMP     : real := 5000.0;  -- Fixed typo (was 50000.0)
    constant NOISE_FLOOR      : real := 20.0;

    -- =========================================================================
    -- Signals
    -- =========================================================================
    signal aclk    : std_logic := '0';
    signal aresetn : std_logic := '0';
    
    signal s_axis_tdata  : std_logic_vector(31 downto 0) := (others => '0');
    signal s_axis_tvalid : std_logic := '0';
    signal s_axis_tlast  : std_logic := '0';
    signal s_axis_tready : std_logic;
    
    signal m_axis_tdata    : std_logic_vector(16 downto 0);
    signal m_axis_tvalid   : std_logic;
    signal m_axis_tlast    : std_logic;
    signal m_axis_tready   : std_logic := '1';
    
    signal rdm_range_bin   : std_logic_vector(9 downto 0);
    signal rdm_doppler_bin : std_logic_vector(6 downto 0);
    
    signal status_range_fft_done   : std_logic;
    signal status_doppler_fft_done : std_logic;
    signal status_frame_complete   : std_logic;
    signal status_overflow         : std_logic;
    
    signal sim_done : std_logic := '0';
    signal output_sample_count : integer := 0;

    -- Timeout watchdog
    constant TIMEOUT_CYCLES : integer := 10000000;  -- 100ms at 100MHz

begin

    -- =========================================================================
    -- DUT Instantiation
    -- =========================================================================
    uut: radar_core_v3
    generic map (
        N_RANGE   => N_RANGE,
        N_DOPPLER => N_DOPPLER
    )
    port map (
        aclk            => aclk,
        aresetn         => aresetn,
        s_axis_tdata    => s_axis_tdata,
        s_axis_tvalid   => s_axis_tvalid,
        s_axis_tlast    => s_axis_tlast,
        s_axis_tready   => s_axis_tready,
        m_axis_tdata    => m_axis_tdata,
        m_axis_tvalid   => m_axis_tvalid,
        m_axis_tlast    => m_axis_tlast,
        m_axis_tready   => m_axis_tready,
        rdm_range_bin   => rdm_range_bin,
        rdm_doppler_bin => rdm_doppler_bin,
        status_range_fft_done   => status_range_fft_done,
        status_doppler_fft_done => status_doppler_fft_done,
        status_frame_complete   => status_frame_complete,
        status_overflow         => status_overflow
    );

    -- =========================================================================
    -- Clock Generation
    -- =========================================================================
    clk_proc: process
    begin
        while sim_done = '0' loop
            aclk <= '0';
            wait for CLK_PERIOD/2;
            aclk <= '1';
            wait for CLK_PERIOD/2;
        end loop;
        wait;
    end process;

    -- =========================================================================
    -- Stimulus Process - GATED (no magic waits)
    -- =========================================================================
    stimulus_proc: process
        variable seed1, seed2 : positive := 1;
        variable rand : real;
        variable chirp_num : integer;
        variable sample_num : integer;
        variable i_acc, q_acc : real;
        variable phase : real;
        variable i_val, q_val : integer;
    begin
        -- Reset sequence
        aresetn <= '0';
        s_axis_tvalid <= '0';
        s_axis_tlast <= '0';
        
        -- Wait for clock to stabilize (sync to edge, not time-based)
        wait until rising_edge(aclk);
        wait until rising_edge(aclk);
        wait until rising_edge(aclk);
        
        aresetn <= '1';
        
        -- GATED: Wait for core to indicate readiness via tready
        -- This replaces magic time-based waits
        report "Waiting for core readiness (s_axis_tready = '1')...";
        wait until s_axis_tready = '1' and rising_edge(aclk);
        
        report "Core ready. Starting data transmission.";
        
        -- Generate 1 CPI for testing (change to 2 for full test)
        for cpi in 0 to 0 loop
            report "=== Generating CPI " & integer'image(cpi) & " ===";
            
            for chirp_num in 0 to N_DOPPLER-1 loop
                for sample_num in 0 to N_RANGE-1 loop
                    i_acc := 0.0;
                    q_acc := 0.0;
                    
                    -- Target 1
                    phase := 2.0 * MATH_PI * (
                        real(TARGET_1_RANGE) * real(sample_num) / real(N_RANGE) +
                        TARGET_1_DOPPLER * real(chirp_num) / real(N_DOPPLER)
                    );
                    i_acc := i_acc + TARGET_1_AMP * cos(phase);
                    q_acc := q_acc + TARGET_1_AMP * sin(phase);
                    
                    -- Target 2
                    phase := 2.0 * MATH_PI * (
                        real(TARGET_2_RANGE) * real(sample_num) / real(N_RANGE) +
                        TARGET_2_DOPPLER * real(chirp_num) / real(N_DOPPLER)
                    );
                    i_acc := i_acc + TARGET_2_AMP * cos(phase);
                    q_acc := q_acc + TARGET_2_AMP * sin(phase);
                    
                    -- Noise
                    uniform(seed1, seed2, rand);
                    i_acc := i_acc + NOISE_FLOOR * (rand - 0.5) * 2.0;
                    uniform(seed1, seed2, rand);
                    q_acc := q_acc + NOISE_FLOOR * (rand - 0.5) * 2.0;
                    
                    -- Quantize and clamp
                    i_val := integer(i_acc);
                    q_val := integer(q_acc);
                    if i_val > 32767 then i_val := 32767; elsif i_val < -32768 then i_val := -32768; end if;
                    if q_val > 32767 then q_val := 32767; elsif q_val < -32768 then q_val := -32768; end if;
                    
                    -- Drive AXI-Stream with proper handshaking
                    s_axis_tdata <= std_logic_vector(to_signed(q_val, 16)) & std_logic_vector(to_signed(i_val, 16));
                    s_axis_tvalid <= '1';
                    s_axis_tlast <= '1' when sample_num = N_RANGE-1 else '0';
                    
                    -- GATED handshake: wait for ready
                    wait until rising_edge(aclk);
                    while s_axis_tready = '0' loop
                        wait until rising_edge(aclk);
                    end loop;
                end loop;
            end loop;
        end loop;
        
        s_axis_tvalid <= '0';
        s_axis_tlast <= '0';
        
        report "Data transmission complete. Waiting for processing...";
        
        -- GATED: Wait for frame complete signal (not time-based)
        wait until status_frame_complete = '1' and rising_edge(aclk);
        
        -- Allow output pipeline to drain
        for i in 0 to 1000 loop
            wait until rising_edge(aclk);
            exit when m_axis_tvalid = '0';
        end loop;
        
        sim_done <= '1';
        report "===== Simulation Complete =====";
        report "Total output samples: " & integer'image(output_sample_count);
        if status_overflow = '1' then
            report "WARNING: Overflow detected in pipeline!" severity warning;
        else
            report "No overflow detected - bit growth managed correctly.";
        end if;
        wait;
    end process;

    -- =========================================================================
    -- Timeout Watchdog
    -- =========================================================================
    watchdog_proc: process
        variable cycle_count : integer := 0;
    begin
        wait until aresetn = '1';
        while sim_done = '0' loop
            wait until rising_edge(aclk);
            cycle_count := cycle_count + 1;
            if cycle_count > TIMEOUT_CYCLES then
                report "TIMEOUT: Simulation exceeded maximum cycles" severity failure;
            end if;
        end loop;
        wait;
    end process;

    -- =========================================================================
    -- Output Monitor
    -- =========================================================================
    monitor_proc: process
        file output_file : text open write_mode is "radar_output.txt";
        variable outline : line;
        variable mag_val : integer;
        variable range_idx : integer;
        variable doppler_idx : integer;
    begin
        wait until aresetn = '1';
        
        loop
            wait until rising_edge(aclk);
            exit when sim_done = '1';
            
            if m_axis_tvalid = '1' and m_axis_tready = '1' then
                mag_val := to_integer(unsigned(m_axis_tdata));
                range_idx := to_integer(unsigned(rdm_range_bin));
                doppler_idx := to_integer(unsigned(rdm_doppler_bin));
                
                write(outline, range_idx);
                write(outline, string'(" "));
                write(outline, doppler_idx);
                write(outline, string'(" "));
                write(outline, mag_val);
                writeline(output_file, outline);
                
                output_sample_count <= output_sample_count + 1;
                
                if mag_val > 50000 then
                     report "Target Detected! R=" & integer'image(range_idx) & 
                            " D=" & integer'image(doppler_idx) & 
                            " Mag=" & integer'image(mag_val);
                end if;
            end if;
        end loop;
        
        file_close(output_file);
        wait;
    end process;

end Behavioral;